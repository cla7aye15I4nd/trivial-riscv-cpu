module cpu_if(
    input wire clk,
    input wire rdy,
    input wire rst,
    
    input wire hitx,
    input wire hity,
    input wire `word_t instx,
    input wire `word_t insty,

    output wire en_rx_out,
    output wire en_ry_out,
    output wire `addr_t pcx_out,
    output wire `addr_t pcy_out,

    output reg `inst_t pc0_out,
    output reg `inst_t pc1_out,
    output reg hitx_out,
    output reg hity_out,
    output reg `word_t instx_out,
    output reg `word_t insty_out
);

reg `addr_t pcx, pcy;

assign en_rx_out = 1;
assign en_ry_out = 1;
assign pcx_out = pcx;
assign pcy_out = pcy;

`define REV(inst) {inst[7 : 0], inst[15 : 8], inst[23: 16], inst[31 : 24]}
always @(posedge clk) begin
    if (rst) begin
        pcx <= 0;
        pcy <= 4;
    end else if (rdy) begin
        pc0_out <= pcx;
        pc1_out <= pcy;
        if (hitx) begin
            hitx_out  <= 1;
            instx_out <= `REV(instx);
            if (hity) begin
                hity_out  <= 1;
                insty_out <= `REV(insty);
                pcx <= pcx + 8;
                pcy <= pcy + 8;
            end else begin
                hity_out  <= 0;
                insty_out <= `ZERO_WORD;
                pcx <= pcx + 4;
                pcy <= pcy + 4;
            end
        end else begin
            instx_out <= `ZERO_WORD;
            hitx_out <= 0;
            hity_out <= 0;
        end
    end
end
endmodule // cpu_if